module Regfile (
    ports
);
    
endmodule