`include "defines.v"
module ex_stage (
    
);
    
endmodule