

module cache{
   input write_addr,
   input read_addr,
   input write_en,
   input read_en,
   input write_data,
   output read_data, 
   input write_mask,

   output axi_write_addr,
   output axi_read_addr,
   output axi_
   
}